.title KiCad schematic
M4 Net-_M1-Pad1_ /B /VDD /VDD PMOS_OR1 l=1u w=6u
M1 Net-_M1-Pad1_ /A /VDD /VDD PMOS_OR1 l=1u w=6u
M2 Net-_M1-Pad1_ /A /X /X NMOS_OR1 l=1u w=2u
M3 /X /B /VSS /VSS NMOS_OR1 l=1u w=2u
.end
